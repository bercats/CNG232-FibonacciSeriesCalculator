library verilog;
use verilog.vl_types.all;
entity FSM_DECO_tb is
end FSM_DECO_tb;
