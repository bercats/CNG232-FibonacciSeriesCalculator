library verilog;
use verilog.vl_types.all;
entity FSM_tb is
end FSM_tb;
