library verilog;
use verilog.vl_types.all;
entity FIBO_FSM_tb is
end FIBO_FSM_tb;
