library verilog;
use verilog.vl_types.all;
entity decoder_2to4_tb is
end decoder_2to4_tb;
