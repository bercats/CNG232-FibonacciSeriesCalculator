library verilog;
use verilog.vl_types.all;
entity mux_2to1_tb is
end mux_2to1_tb;
